// Can be adjusted, but the array size below needs to be the same number
const int CAP = 100;

f<int> main() {
    int[CAP] board;

    // Initialize board
    for int i = 0; i < CAP; i++ {
        board[i] = 0;
    }
    board[CAP - 2] = 1; // Set second-last element to 1

    // Print pattern
    for int i = 0; i < CAP - 2; i++ {
        for int j = 0; j < CAP; j++ {
            printf("%s", board[j] == 1 ? "*" : " ");
        }
        printf("\n");

        int pattern = (board[0] << 1) | board[1];
        for int j = 1; j < CAP - 1; j++ {
            pattern = ((pattern << 1) & 7) | board[j + 1];
            board[j] = (110 >> pattern) & 1;
        }
    }
}
// Inspired by: https://www.geeksforgeeks.org/program-for-conways-game-of-life

import "std/math/rand" as rand;

const int row = 10;
const int col = 10;
const int generationsToCalculate = 5;

p rowLineTop() {
    printf("\n");
    for int i = 0; i < col; i++ { printf("╭─────╮"); }
    printf("\n");
}

p rowLineMiddle() {
    printf("\n");
    for int i = 0; i < col; i++ { printf("├─────┤"); }
    printf("\n");
}

p rowLineBottom() {
    printf("\n");
    for int i = 0; i < col; i++ { printf("╰─────╯"); }
    printf("\n");
}

p printGeneration(string name, int[10][10] matrix) {
    printf("%s:\n", name);
    rowLineTop();
    for int i = 0; i < row; i++ {
        if i > 0 {
            rowLineMiddle();
        }
        for int j = 0; j < col; j++ {
            printf("│  %d  │", matrix[i][j]);
        }
    }
    rowLineBottom();
}

f<int> countLiveNeighborCell(int[10][10] matrix, int r, int c) {
    int count = 0;
    for int i = r - 1; i <= r + 1; i++ {
        for int j = c - 1; j <= c + 1; j++ {
            if (i == r && j == c) || (i < 0 || j < 0) || (i >= row || j >= col) {
                continue;
            }
            if matrix[i][j] == 1 {
                count++;
            }
        }
    }
    return count;
}

f<int> main() {
    int[10][10] a;
    int[10][10] b;

    // Generate matrix canvas with random values (live and dead cells)
    for int i = 0; i < row; i++ {
        for int j = 0; j < col; j++ {
            a[i][j] = rand.randInt(0, 1);
        }
    }
    printGeneration("Initial state", a);

    for int generation = 1; generation < generationsToCalculate; generation++ {
        // Calculate next generation
        for int i = 0; i < row; i++ {
            for int j = 0; j < col; j++ {
                int neighbor_live_cell = countLiveNeighborCell(a, i, j);
                if a[i][j] == 1 && (neighbor_live_cell == 2 || neighbor_live_cell == 3) {
                    b[i][j] = 1;
                } else if a[i][j] == 0 && neighbor_live_cell == 3 {
                    b[i][j] = 1;
                } else {
                    b[i][j] = 0;
                }
            }
        }

        // Print next generation
        printGeneration("\nNext generation", b);

        // Set new matrix to old matrix
        a = b;
    }
}

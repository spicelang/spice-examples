// Inspired by GeeksForGeeks: https://www.geeksforgeeks.org/sudoku-backtracking-7

const int size = 9;

p print(int[][] grid) {
    for int i = 0; i < size; i++ {
        for int j = 0; j < size; j++ {
             printf("%d ", grid[i][j]);
        }
        printf("\n");
    }
}

f<bool> isSafe(int[][] grid, int row, int col, int num) {
    // Check if we find the same num in the similar row -> return false
    for int x = 0; x <= size - 1; x++ {
        if grid[row][x] == num {
            return false;
        }
    }

    // Check if we find the same num in the similar column -> return false
    for int x = 0; x <= size - 1; x++ {
        if grid[x][col] == num {
            return false;
        }
    }

    // Check if we find the same num in the particular 3*3 matrix -> return false
    int startRow = row - row % 3;
    int startCol = col - col % 3;

    for int i = 0; i < 3; i++ {
        for int j = 0; j < 3; j++ {
            if grid[i + startRow][j + startCol] == num {
                return false;
            }
        }
    }

    return true;
}

f<bool> solveSudoku(int[][] grid, int row, int col) {
    // Check if we have reached the second last row and the last column.
    // We return true to avoid further backtracking
    if row == size - 1 && col == size { return true; }

    if col == size {
        row++;
        col = 0;
    }

    if grid[row][col] > 0 {
        return solveSudoku(grid, row, col + 1);
    }

    for int num = 1; num <= size; num++ {
        if isSafe(grid, row, col, num) {
            grid[row][col] = num;

            if solveSudoku(grid, row, col + 1) {
                return true;
            }
        }
        grid[row][col] = 0;
    }

    return false;
}

f<int> main() {
    int[size][size] grid = {
        { 3, 0, 6, 5, 0, 8, 4, 0, 0 },
        { 5, 2, 0, 0, 0, 0, 0, 0, 0 },
        { 0, 8, 7, 0, 0, 0, 0, 3, 1 },
        { 0, 0, 3, 0, 1, 0, 0, 8, 0 },
        { 9, 0, 0, 8, 6, 3, 0, 0, 5 },
        { 0, 5, 0, 0, 9, 0, 6, 0, 0 },
        { 1, 3, 0, 0, 0, 0, 2, 5, 0 },
        { 0, 0, 0, 0, 0, 0, 0, 7, 4 },
        { 0, 0, 5, 2, 0, 6, 3, 0, 0 }
    };

    if solveSudoku(grid, 0, 0) {
        print(grid);
    } else {
        printf("No solution was found.");
    }
}